Require Export Protocol.
Require Export Uint63.
Require Extraction.
Extraction Blacklist Uint63 List String.

Include Protocol.

Require ExtrOcamlBasic.
Require ExtrOcamlNativeString.
Require ExtrOCamlInt63.
Require ExtrOcamlZInt.

(* This is necessary to do proper extraction of the Coq representation
   of the file_descr Unix type. *)
Extract Constant ProtocolDefinitions.file_descr => "Unix.file_descr".
Extract Constant ProtocolDefinitions.sockaddr => "Unix.sockaddr".
Extract Constant ProtocolDefinitions.eqb_sockaddr => "fun x y -> x = y".


(*Extract Constant Uint63.Uint63.t => "int".*)


(*
Extraction Library ProtocolDefinitions.
 *)

(* To avoid errors like


File "Protocol.mli", line 1, characters 5-14:
1 | open Datatypes
         ^^^^^^^^^
Error: Unbound module Datatypes


we have to provide access to Datatypes module. This module
can be automatically generated by Coq extraction, but
we have to trigger its recursive version. *)
Recursive Extraction Library Protocol.

(* 
This must be accompanied by a scheme that properly establishes
the compilation dependencies for the generated files. Therefore
we added the depend target to Makefile.

We also have to add many more items to clean.
*)


(*
This is done now by the library extraction:
Recursive Extraction dir_to_string. *)
